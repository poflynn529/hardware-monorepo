package utils;

function automatic int cdiv(int numerator, int denominator);
    return (numerator + denominator - 1) / denominator;
endfunction

endpackage
